library verilog;
use verilog.vl_types.all;
entity testebench_somador is
end testebench_somador;

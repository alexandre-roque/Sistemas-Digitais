library verilog;
use verilog.vl_types.all;
entity testebench_registrador is
end testebench_registrador;
